module mirror_spi_driver(clk, ss, datain, dataout);











endmodule 