module Font_library(VGA_clk, currentLetter, xPixel, yPixel, pixelOutput);
	input VGA_clk;
	input [6:0] currentLetter;
	input [9:0] xPixel, yPixel;
	
	output pixelOutput;
	
	wire [0:40447]font_library;
	
	initialize_fonts(font_library);
	
	assign pixelOutput = font_library[{currentLetter, yPixel[4:0], xPixel[3:0]}];

endmodule


//[^\d]+
//http://ece320web.groups.et.byu.net/labs/VGATextGeneration/list_ch13_01_font_rom.vhd
module initialize_fonts(font_library);

	output [0:40447] font_library;
	assign font_library = 40448'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000001111000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000011000000000000111100000000000011110000000000111100000000000011110000000000111100000000000011110000000000111100000000000011110000000000111100000000000011110000000000111100000000000011110000000000001100000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110000111100000011110011110000001111001111000000111100111100000011110011110000111111001111000011111100111100111111110011110011111111001111111100111100111111110011110011111100001111001111110000111100111100000011110011110000001111001111000000111100111100000011110000111111111100000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000011110000000000111111000000000011111100000000111111110000000011111111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000001111111111110000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000001111111111000011110000001111001111000000111100000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000000111100000011110011110000001111001111111111111100111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110000111100000011110011110000001111000000000000111100000000000011110000000000001111000000000000111100000011111111000000001111111100000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111001111000000111100111100000011110000111111111100000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000111100000000001111110000000000111111000000001111111100000000111111110000001111001111000000111100111100001111000011110000111100001111000011111111111111001111111111111100000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000111111110000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100111111111111110011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011111111111100001111111111110000000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100111100000011110011110000001111000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000111111000000001111000000000000111100000000001111000000000000111100000000000011110000000000001111000000000000111111111111000011111111111100001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110000111111111100000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110011111111111111001111000000111100111100000011110000000000001111000000000000111100000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000001111111111000011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110000111111111100000011111111110000111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110000111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100001111111111110000111111111111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000011110000000000001111000000111111110000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000111100000000000011110000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000011110000000000001111000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000111100000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000000001111000000000000111100000000000000111100000000000011110000000000000011110000000000001111000000000000001111000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000111111111111000000000000000000000000000000000000000000000000000000000000000000001111111111110000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000011110000000000000011110000000000001111000000000000001111000000000000111100000000000000111100000000000011110000000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110000111100000011110011110000001111001111000000111100111100000011110000000000111100000000000011110000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000000000000000000000000000000000001111000000000000111100000000000011110000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000111111111100001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111001111111100111100111111110011110011111111001111001111111100111100111111110011110011111111001111001111110000111100111111000011110000000000001111000000000000001111111111000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000110000000000001111110000000000111111000000001111001111000000111100111100001111000000111100111100000011110011110000001111001111000000111100111111111111110011111111111111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100001111111111110000001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111111111000000111111111100000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110011111111111100001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001111111100000011110000111100001111000011110011110000000011001111000000001100111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000001100111100000000110000111100001111000011110000111100000011111111000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000111111111100000000111100111100000011110011110000001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111001111000000111100111100001111111111000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111111111100001111000011110000111100001111000011110000001100001111000000110000111100110000000011110011000000001111111100000000111111110000000011110011000000001111001100000000111100000000000011110000000000001111000000110000111100000011000011110000111100001111000011110011111111111111001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110011111111111111000011110000111100001111000011110000111100000011000011110000001100001111001100000000111100110000000011111111000000001111111100000000111100110000000011110011000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000111111110000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000011111111000000111100001111000011110000111100111100000000110011110000000011001111000000000000111100000000000011110000000000001111000000000000111100111111110011110011111111001111000000111100111100000011110011110000001111001111000000111100001111000011110000111100001111000000111111001100000011111100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111111111111110011111111111111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001111111100000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000011111111000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000111111110000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100000011111111000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100001111001111110000111100001111000011110000111100001111000011110000111100001111000011110000111100111100000011110011110000001111111100000000111111110000000011111111000000001111111100000000111100111100000011110011110000001111000011110000111100001111000011110000111100001111000011110011111100001111001111110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000011111111000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000001100001111000000110000111100001111000011110000111100111111111111110011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000011100111000000001110011110000001111001111100001111100111110000111110011111100111111001111111111111100111111111111110011111111111111001110011110011100111001111001110011100011000111001110000000011100111000000001110011100000000111001110000000011100111000000001110011100000000111001110000000011100111000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000001111001111000000111100111111000011110011111100001111001111111100111100111111110011110011111111111111001111111111111100111100111111110011110011111111001111000011111100111100001111110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000111111111100001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100001111111111000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000111111111111000000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111111111100000011111111110000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000001111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110000111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100110011110011110011001111001111001111111100111100111111110000111111111100000011111111110000000000001111000000000000111100000000000011111100000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000011111111111100000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011111111110000001111111111000000111100111100000011110011110000001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100111111000011110011111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000001111111111000011110000001111001111000000111100111100000011110011110000001111000011110000000000001111000000000000001111110000000000111111000000000000001111000000000000111100000000000000111100000000000011110011110000001111001111000000111100111100000011110011110000001111000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111111111100111111111111110011100111100111001110011110011100000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000011111111000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100001111111111000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000011100111000000001110011100000000111001110000000011100111000000001110011100000000111001110000000011100111000000001110011100000000111001110000000011100111000000001110011100000000111001110000000011100111000000001110001110000001110000111100001111000000111001110000000011111111000000000011110000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000111001110000000011100111000000001110011100000000111001110000000011100111000000001110011100000000111001110000000011100111000000001110011100000000111001110001100011100111001111001110011100111100111001110011110011100111111111111110011111100111111000111100001111000011110000111100001111000011110000111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000001110011100000000111001110000000011100111000000001110001111000011110000111100001111000000111111110000000011111111000000000011110000000000001111000000000000111100000000000011110000000000111111110000000011111111000000111100001111000011110000111100011100000000111001110000000011100111000000001110011100000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000011100111000000001110011100000000111001110000000011100111000000001110011100000000111000111100001111000011110000111100000011100111000000001111111100000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000001111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111111111100111000000001110011100000000111001000000001111000000000000111100000000001111000000000000111100000000001111000000000000111100000000001111000000000000111100000000001111000000000000111100000000000111000000000000011100000000001001110000000011100111000000001110011111111111111001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001111111100000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011111111000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000001100000000000000111100000000000011110000000000001111110000000000111111000000000000111111000000000011111100000000000011111100000000001111110000000000001111110000000000111111000000000000111111000000000011111100000000000011110000000000001111000000000000001100000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000111111110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000001111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000110000000000001111110000000000111111000000001111001111000000111100111100001111000000111100111100000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000000011110000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000111111110000000000000011110000000000001111000000111111111100000011111111110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000001111110011110000111111001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000111111000000000000111100000000000011110000000000001111000000000000111100000000000011111111000000001111111100000000111100111100000011110011110000001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110000111100000011110011110000001111001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000111100111100000011110000111111111100000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000011111100000000000011110000000000001111000000000000111100000000000011110000000011111111000000001111111100000011110011110000001111001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000001111110011110000111111001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000001111111111000011110000001111001111000000111100111111111111110011111111111111001111000000000000111100000000000011110000000000001111000000000000111100000011110011110000001111000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000111111000000001111001111000000111100111100000011110000110000001111000011000000111100000000000011110000000000111111110000000011111111000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000011111111000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110011110000111111001111001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000001111111111000000111111111100000000000011110000000000001111000011110000111100001111000011110000001111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000111111000000000000111100000000000011110000000000001111000000000000111100000000000011110011110000001111001111000000111111001111000011111100111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111001111110000111100111111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000001111110000000000111111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000001111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000001111110000000000111111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000011110000111100001111000011110000111100001111000011110000111100000011111111000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000111111000000000000111100000000000011110000000000001111000000000000111100000000000011110000111100001111000011110000111100111100000011110011110000001111111100000000111111110000000011111111000000001111111100000000111100111100000011110011110000001111000011110000111100001111001111110000111100111111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000111111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000001111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000011110011111100001111001111111111111111111111111111111111110011110011111111001111001111111100111100111111110011110011111111001111001111111100111100111111110011110011111111001111001111111100111100111111110011110011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111001111110000111100111111000000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000011111111110000111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110000111111111100000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100111111000011110011111100000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111111111000000111111111100000011110000000000001111000000000000111100000000000011110000000000111111110000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100111100001111110011110011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100000011111111110000001111111111000000000000111100000000000011110000000000001111000000000000111100000000001111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110011111100001111001111110000001111110011110000111111001111000011110000111100001111000011110000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000011111111000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000111111111100001111000000111100111100000011110000111100000000000011110000000000000011111100000000001111110000000000000011110000000000001111000011110000001111001111000000111100001111111111000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000110000000000001111000000000000111100000000000011110000000000001111000000001111111111110000111111111111000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110011110000001111001111000000001111110000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000000111111001111000011111100111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000111111110000000011111111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011110011110000111100001111000011110000001111111100000000111111110000000000111100000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000001111111100000000111111110000000011111111000000001111111100000000111111110000000011111111001111001111111100111100111111110011110011111111001111001111111111111111111111111111111111110011110000111100001111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000011111111000000001111001111000011110000111100001111000000111111110000000011111111000000000011110000000000001111000000000011111111000000001111111100000011110000111100001111000011110011110000000011111111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100001111111111110000111111111111000000000000111100000000000011110000000000111100000000000011110000111111111100000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100111111111111110011110000111100001111000011110000000000111100000000000011110000000000111100000000000011110000000000111100000000000011110000000000111100000011110011110000001111001111111111111100111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//	//0 = 000000
//	assign font_library[0:511] = 512'b00000000000000000000000000000000000000000000000000000000000000000011111111110000001111111111000011110000001111001111000000111100111100000011110011110000001111001111000011111100111100001111110011110011111111001111001111111100111111110011110011111111001111001111110000111100111111000011110011110000001111001111000000111100111100000011110011110000001111000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//	
//	//1 = 000001
//	assign font_library[512:1023] = 512'b00000000000000000000000000000000000000000000000000000000000000000000001111000000000000111100000000001111110000000000111111000000001111111100000000111111110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000011111111111100001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//	
//	//2 = 000010
//	assign font_library[1024:1535] = 512'b00000000000000000000000000000000000000000000000000000000000000000011111111110000001111111111000011110000001111001111000000111100000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000000111100000011110011110000001111001111111111111100111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//
//	//3 = 000011
//	assign font_library[1536:2047] = 512'b00000000000000000000000000000000000000000000000000000000000000000011111111110000001111111111000011110000001111001111000000111100000000000011110000000000001111000000000000111100000000000011110000001111111100000000111111110000000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100111100000011110011110000001111000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//	
//	//4 = 000100
//	assign font_library[2048:2559] = 512'b00000000000000000000000000000000000000000000000000000000000000000000000011110000000000001111000000000011111100000000001111110000000011111111000000001111111100000011110011110000001111001111000011110000111100001111000011110000111100001111110011111111111111001111111111111100000000001111000000000000111100000000000011110000000000001111000000000000111100000000001111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//	
//	//5 = 000101
//	assign font_library[2560:3071] = 512'b00000000000000000000000000000000000000000000000000000000000000001111111111111100111111111111110011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011111111111100001111111111110000000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100111100000011110011110000001111000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//	
//	//6 = 000110
//	assign font_library[3072:3583] = 512'b00000000000000000000000000000000000000000000000000000000000000000000111111000000000011111100000000111100000000000011110000000000111100000000000011110000000000001111000000000000111100000000000011111111111100001111111111110000111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//	
//	//7 = 000111
//	assign font_library[3584:4095] = 512'b00000000000000000000000000000000000000000000000000000000000000001111111111111100111111111111110011110000001111001111000000111100000000000011110000000000001111000000000000111100000000000011110000000000111100000000000011110000000000111100000000000011110000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//	
//	//8 = 001000
//	assign font_library[4096:4607] = 512'b00000000000000000000000000000000000000000000000000000000000000000011111111110000001111111111000011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110000111111111100000011111111110000111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110011110000001111000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//	
//	//9 = 001001
//	assign font_library[4608:5119] = 512'b00000000000000000000000000000000000000000000000000000000000000000011111111110000001111111111000011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110000111111111110000011111111111000000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000001111000000000000111100000011111111000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//	
//	//A = 001010
//	assign font_library[5120:5631] = 512'b00000000000000000000000000000000000000000000000000000000000000000000001100000000000001111000000000001111110000000000111111000000001111001111000000111100111100001111000000111100111100000011110011110000001111001111000000111100111100000011110011111111111111001111111111111100111100000011110011110000001111001111000000111100111100000011110011110000001111001111000000111100111100000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//	
//	//B = 001011
//	assign font_library[5632:6143] = 512'b00000000000000000000000000000000000000000000000000000000000000001111111111110000111111111111000000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111111111100000011111111110000001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111001111111111110000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//	
//	//C = 001100
//	assign font_library[6144:6655] = 512'b00000000000000000000000000000000000000000000000000000000000000000000111111110000000011111111000000111100001111000011110000111100111100000000110011110000000011001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000011001111000000001100001111000011110000111100001111000000111111110000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//
//	//D = 001101
//	assign font_library[6656:7167] = 512'b00000000000000000000000000000000000000000000000000000000000000001111111111000000111111111100000000111100111100000011110011110000001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111000011110000111100001111101111000000111110111100001111111111000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//	
//	//E = 001110
//	assign font_library[7168:7679] = 512'b00000000000000000000000000000000000000000000000000000000000000001111111111111100111111111111110000111100001111000011110000111100001111000000110000111100000011000011110011000000001111001100000000111111110000000011111111000000001111001100000000111100110000000011110000000000001111000000000000111100000011000011110000001100001111000011110000111100001111001111111111111100111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//	
//	//F = 001111
//	assign font_library[7680:8191] = 512'b00000000000000000000000000000000000000000000000000000000000000001111111111111100111111111111110000111100001111000011110000111100001111000000110000111100000011000011110011000000001111001100000000111111110000000011111111000000001111001100000000111100110000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000001111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//	
	endmodule
