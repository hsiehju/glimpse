module Font_library(VGA_clk, currentLetter, xPixel, yPixel, pixelOutput);
	input VGA_clk;
	input [5:0] currentLetter;
	input [9:0] xPixel, yPixel;
	
	output pixelOutput;
	
	wire [0:20991]font_library;
	
	initialize_fonts(font_library);
	
	assign pixelOutput = font_library[{currentLetter, yPixel[4:0], xPixel[3:0]}];

endmodule


//[^\d]+
//http://ece320web.groups.et.byu.net/labs/VGATextGeneration/list_ch13_01_font_rom.vhd
module initialize_fonts(font_library);

	output [0:20991] font_library;
	//0 = 000000
	assign font_library[0:511] = 512'b00000000000000000000000000000000000000000000000000000000000000000011111111110000001111111111000011110000001111001111000000111100111100000011110011110000001111001111000011111100111100001111110011110011111111001111001111111100111111110011110011111111001111001111110000111100111111000011110011110000001111001111000000111100111100000011110011110000001111000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	//1 = 000001
	assign font_library[512:1023] = 512'b00000000000000000000000000000000000000000000000000000000000000000000001111000000000000111100000000001111110000000000111111000000001111111100000000111111110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000011111111111100001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	//2 = 000010
	assign font_library[1024:1535] = 512'b00000000000000000000000000000000000000000000000000000000000000000011111111110000001111111111000011110000001111001111000000111100000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000011110000000000001111000000000000111100000011110011110000001111001111111111111100111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

	//3 = 000011
	assign font_library[1536:2047] = 512'b00000000000000000000000000000000000000000000000000000000000000000011111111110000001111111111000011110000001111001111000000111100000000000011110000000000001111000000000000111100000000000011110000001111111100000000111111110000000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100111100000011110011110000001111000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	//4 = 000100
	assign font_library[2048:2559] = 512'b00000000000000000000000000000000000000000000000000000000000000000000000011110000000000001111000000000011111100000000001111110000000011111111000000001111111100000011110011110000001111001111000011110000111100001111000011110000111100001111110011111111111111001111111111111100000000001111000000000000111100000000000011110000000000001111000000000000111100000000001111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	//5 = 000101
	assign font_library[2560:3071] = 512'b00000000000000000000000000000000000000000000000000000000000000001111111111111100111111111111110011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000011111111111100001111111111110000000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100111100000011110011110000001111000011111111110000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
endmodule
